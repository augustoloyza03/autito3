library verilog;
use verilog.vl_types.all;
entity SumaoResta_vlg_vec_tst is
end SumaoResta_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ubicacionparte2_vlg_check_tst is
    port(
        SorR            : in     vl_logic;
        Z0              : in     vl_logic;
        Z1              : in     vl_logic;
        Z2              : in     vl_logic;
        Z3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ubicacionparte2_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity ubicacionparte2_vlg_vec_tst is
end ubicacionparte2_vlg_vec_tst;

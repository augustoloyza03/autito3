library verilog;
use verilog.vl_types.all;
entity pruebaadc_vlg_vec_tst is
end pruebaadc_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ubicacionparte2v2_vlg_vec_tst is
end ubicacionparte2v2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity doblar2_vlg_vec_tst is
end doblar2_vlg_vec_tst;

-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sat Nov 09 22:14:14 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ubicacionparte2 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Gizq : IN STD_LOGIC := '0';
        Gder : IN STD_LOGIC := '0';
        S : IN STD_LOGIC := '0';
        Z3 : OUT STD_LOGIC;
        Z2 : OUT STD_LOGIC;
        Z1 : OUT STD_LOGIC;
        Z0 : OUT STD_LOGIC;
        SorR : OUT STD_LOGIC
    );
END ubicacionparte2;

ARCHITECTURE BEHAVIOR OF ubicacionparte2 IS
    TYPE type_fstate IS (O1,O2,O3,O4,RESTAR1,SUMAR4,SUMAR1,RESTAR4);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Gizq,Gder,S)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= O1;
            Z3 <= '0';
            Z2 <= '0';
            Z1 <= '0';
            Z0 <= '0';
            SorR <= '0';
        ELSE
            Z3 <= '0';
            Z2 <= '0';
            Z1 <= '0';
            Z0 <= '0';
            SorR <= '0';
            CASE fstate IS
                WHEN O1 =>
                    IF ((S = '1')) THEN
                        reg_fstate <= O1;
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR1;
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR4;
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR1;
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= O1;
                    END IF;

                    IF ((S = '1')) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((S = '1')) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN O2 =>
                    IF ((S = '1')) THEN
                        reg_fstate <= O2;
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR1;
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR4;
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR1;
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= O2;
                    END IF;

                    IF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    ELSIF ((S = '1')) THEN
                        Z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((S = '1')) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN O3 =>
                    IF ((S = '1')) THEN
                        reg_fstate <= O3;
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR1;
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR4;
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR1;
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= O3;
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    ELSIF ((S = '1')) THEN
                        Z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((S = '1')) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN O4 =>
                    IF ((S = '1')) THEN
                        reg_fstate <= O4;
                    ELSIF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR1;
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        reg_fstate <= RESTAR4;
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR1;
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        reg_fstate <= SUMAR4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= O4;
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z2 <= '1';
                    ELSIF ((S = '1')) THEN
                        Z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z1 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        SorR <= '1';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        SorR <= '0';
                    ELSIF ((S = '1')) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '1';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z0 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF ((((Gizq = '1') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '0') AND (Gder = '0')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((((Gizq = '1') AND (Gder = '1')) AND (S = '0'))) THEN
                        Z3 <= '0';
                    ELSIF ((S = '1')) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN RESTAR1 =>
                    IF ((S = '0')) THEN
                        reg_fstate <= RESTAR1;
                    ELSIF ((S = '1')) THEN
                        reg_fstate <= O2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= RESTAR1;
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN SUMAR4 =>
                    IF ((S = '0')) THEN
                        reg_fstate <= SUMAR4;
                    ELSIF ((S = '1')) THEN
                        reg_fstate <= O1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SUMAR4;
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN SUMAR1 =>
                    IF ((S = '0')) THEN
                        reg_fstate <= SUMAR1;
                    ELSIF ((S = '1')) THEN
                        reg_fstate <= O3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SUMAR1;
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN RESTAR4 =>
                    IF ((S = '0')) THEN
                        reg_fstate <= RESTAR4;
                    ELSIF ((S = '1')) THEN
                        reg_fstate <= O4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= RESTAR4;
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z2 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z1 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        SorR <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        SorR <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z0 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z0 <= '0';
                    END IF;

                    IF (((S = '1') OR (S = '0'))) THEN
                        Z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z3 <= '0';
                    END IF;
                WHEN OTHERS => 
                    Z3 <= 'X';
                    Z2 <= 'X';
                    Z1 <= 'X';
                    Z0 <= 'X';
                    SorR <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;

library verilog;
use verilog.vl_types.all;
entity doblar_vlg_vec_tst is
end doblar_vlg_vec_tst;
